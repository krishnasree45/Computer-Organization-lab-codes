//`include "mux2.v"

module leftbarrelshift32(a,s0,s1,s2,s3,s4,out);

input [31:0]a;
input s0,s1,s2,s3,s4;
output [31:0]out;
wire [31:0]i1,i2,i3,i4;

mux2 ar1(a[31],a[30],s0,i1[31]);
mux2 ar2(a[30],a[29],s0,i1[30]);
mux2 ar3(a[29],a[28],s0,i1[29]);
mux2 ar4(a[28],a[27],s0,i1[28]);
mux2 ar5(a[27],a[26],s0,i1[27]);
mux2 ar6(a[26],a[25],s0,i1[26]);
mux2 ar7(a[25],a[24],s0,i1[25]);
mux2 ar8(a[24],a[23],s0,i1[24]);
mux2 ar9(a[23],a[22],s0,i1[23]);
mux2 ar10(a[22],a[21],s0,i1[22]);
mux2 ar11(a[21],a[20],s0,i1[21]);
mux2 ar12(a[20],a[19],s0,i1[20]);
mux2 ar13(a[19],a[18],s0,i1[19]);
mux2 ar14(a[18],a[17],s0,i1[18]);
mux2 ar15(a[17],a[16],s0,i1[17]);
mux2 ar16(a[16],a[15],s0,i1[16]);
mux2 ar17(a[15],a[14],s0,i1[15]);
mux2 ar18(a[14],a[13],s0,i1[14]);
mux2 ar19(a[13],a[12],s0,i1[13]);
mux2 ar20(a[12],a[11],s0,i1[12]);
mux2 ar21(a[11],a[10],s0,i1[11]);
mux2 ar22(a[10],a[9],s0,i1[10]);
mux2 ar23(a[9],a[8],s0,i1[9]);
mux2 ar24(a[8],a[7],s0,i1[8]);
mux2 ar25(a[7],a[6],s0,i1[7]);
mux2 ar26(a[6],a[5],s0,i1[6]);
mux2 ar27(a[5],a[4],s0,i1[5]);
mux2 ar28(a[4],a[3],s0,i1[4]);
mux2 ar29(a[3],a[2],s0,i1[3]);
mux2 ar30(a[2],a[1],s0,i1[2]);
mux2 ar31(a[1],a[0],s0,i1[1]);
mux2 ar32(a[0],0,s0,i1[0]);




mux2 br1(i1[31],i1[29],s1,i2[31]);
mux2 br2(i1[30],i1[28],s1,i2[30]);
mux2 br3(i1[29],i1[27],s1,i2[29]);
mux2 br4(i1[28],i1[26],s1,i2[28]);
mux2 br5(i1[27],i1[25],s1,i2[27]);
mux2 br6(i1[26],i1[24],s1,i2[26]);
mux2 br7(i1[25],i1[23],s1,i2[25]);
mux2 br8(i1[24],i1[22],s1,i2[24]);
mux2 br9(i1[23],i1[21],s1,i2[23]);
mux2 br10(i1[22],i1[20],s1,i2[22]);
mux2 br11(i1[21],i1[19],s1,i2[21]);
mux2 br12(i1[20],i1[18],s1,i2[20]);
mux2 br13(i1[19],i1[17],s1,i2[19]);
mux2 br14(i1[18],i1[16],s1,i2[18]);
mux2 br15(i1[17],i1[15],s1,i2[17]);
mux2 br16(i1[16],i1[14],s1,i2[16]);
mux2 br17(i1[15],i1[13],s1,i2[15]);
mux2 br18(i1[14],i1[12],s1,i2[14]);
mux2 br19(i1[13],i1[11],s1,i2[13]);
mux2 br20(i1[12],i1[10],s1,i2[12]);
mux2 br21(i1[11],i1[9],s1,i2[11]);
mux2 br22(i1[10],i1[8],s1,i2[10]);
mux2 br23(i1[9],i1[7],s1,i2[9]);
mux2 br24(i1[8],i1[6],s1,i2[8]);
mux2 br25(i1[7],i1[5],s1,i2[7]);
mux2 br26(i1[6],i1[4],s1,i2[6]);
mux2 br27(i1[5],i1[3],s1,i2[5]);
mux2 br28(i1[4],i1[2],s1,i2[4]);
mux2 br29(i1[3],i1[1],s1,i2[3]);
mux2 br30(i1[2],i1[0],s1,i2[2]);
mux2 br31(i1[1],0,s1,i2[1]);
mux2 br32(i1[0],0,s1,i2[0]);

mux2 cr1(i2[31],i2[27],s2,i3[31]);
mux2 cr2(i2[30],i2[26],s2,i3[30]);
mux2 cr3(i2[29],i2[25],s2,i3[29]);
mux2 cr4(i2[28],i2[24],s2,i3[28]);
mux2 cr5(i2[27],i2[23],s2,i3[27]);
mux2 cr6(i2[26],i2[22],s2,i3[26]);
mux2 cr7(i2[25],i2[21],s2,i3[25]);
mux2 cr8(i2[24],i2[20],s2,i3[24]);
mux2 cr9(i2[23],i2[19],s2,i3[23]);
mux2 cr10(i2[22],i2[18],s2,i3[22]);
mux2 cr11(i2[21],i2[17],s2,i3[21]);
mux2 cr12(i2[20],i2[16],s2,i3[20]);
mux2 cr13(i2[19],i2[15],s2,i3[19]);
mux2 cr14(i2[18],i2[14],s2,i3[18]);
mux2 cr15(i2[17],i2[13],s2,i3[17]);
mux2 cr16(i2[16],i2[12],s2,i3[16]);
mux2 cr17(i2[15],i2[11],s2,i3[15]);
mux2 cr18(i2[14],i2[10],s2,i3[14]);
mux2 cr19(i2[13],i2[9],s2,i3[13]);
mux2 cr20(i2[12],i2[8],s2,i3[12]);
mux2 cr21(i2[11],i2[7],s2,i3[11]);
mux2 cr22(i2[10],i2[6],s2,i3[10]);
mux2 cr23(i2[9],i2[5],s2,i3[9]);
mux2 cr24(i2[8],i2[4],s2,i3[8]);
mux2 cr25(i2[7],i2[3],s2,i3[7]);
mux2 cr26(i2[6],i2[2],s2,i3[6]);
mux2 cr27(i2[5],i2[1],s2,i3[5]);
mux2 cr28(i2[4],i2[0],s2,i3[4]);
mux2 cr29(i2[3],0,s2,i3[3]);
mux2 cr30(i2[2],0,s2,i3[2]);
mux2 cr31(i2[1],0,s2,i3[1]);
mux2 cr32(i2[0],0,s2,i3[0]);

mux2 dr1(i3[31],i3[23],s3,i4[31]);
mux2 dr2(i3[30],i3[22],s3,i4[30]);
mux2 dr3(i3[29],i3[21],s3,i4[29]);
mux2 dr4(i3[28],i3[20],s3,i4[28]);
mux2 dr5(i3[27],i3[19],s3,i4[27]);
mux2 dr6(i3[26],i3[18],s3,i4[26]);
mux2 dr7(i3[25],i3[17],s3,i4[25]);
mux2 dr8(i3[24],i3[16],s3,i4[24]);
mux2 dr9(i3[23],i3[15],s3,i4[23]);
mux2 dr10(i3[22],i3[14],s3,i4[22]);
mux2 dr11(i3[21],i3[13],s3,i4[21]);
mux2 dr12(i3[20],i3[12],s3,i4[20]);
mux2 dr13(i3[19],i3[11],s3,i4[19]);
mux2 dr14(i3[18],i3[10],s3,i4[18]);
mux2 dr15(i3[17],i3[9],s3,i4[17]);
mux2 dr16(i3[16],i3[8],s3,i4[16]);
mux2 dr17(i3[15],i3[7],s3,i4[15]);
mux2 dr18(i3[14],i3[6],s3,i4[14]);
mux2 dr19(i3[13],i3[5],s3,i4[13]);
mux2 dr20(i3[12],i3[4],s3,i4[12]);
mux2 dr21(i3[11],i3[3],s3,i4[11]);
mux2 dr22(i3[10],i3[2],s3,i4[10]);
mux2 dr23(i3[9],i3[1],s3,i4[9]);
mux2 dr24(i3[8],i3[0],s3,i4[8]);
mux2 dr25(i3[7],0,s3,i4[7]);
mux2 dr26(i3[6],0,s3,i4[6]);
mux2 dr27(i3[5],0,s3,i4[5]);
mux2 dr28(i3[4],0,s3,i4[4]);
mux2 dr29(i3[3],0,s3,i4[3]);
mux2 dr30(i3[2],0,s3,i4[2]);
mux2 dr31(i3[1],0,s3,i4[1]);
mux2 dr32(i3[0],0,s3,i4[0]);

mux2 er1(i4[31],i4[15],s4,out[31]);
mux2 er2(i4[30],i4[14],s4,out[30]);
mux2 er3(i4[29],i4[13],s4,out[29]);
mux2 er4(i4[28],i4[12],s4,out[28]);
mux2 er5(i4[27],i4[11],s4,out[27]);
mux2 er6(i4[26],i4[10],s4,out[26]);
mux2 er7(i4[25],i4[9],s4,out[25]);
mux2 er8(i4[24],i4[8],s4,out[24]);
mux2 er9(i4[23],i4[7],s4,out[23]);
mux2 er10(i4[22],i4[6],s4,out[22]);
mux2 er11(i4[21],i4[5],s4,out[21]);
mux2 er12(i4[20],i4[4],s4,out[20]);
mux2 er13(i4[19],i4[3],s4,out[19]);
mux2 er14(i4[18],i4[2],s4,out[18]);
mux2 er15(i4[17],i4[1],s4,out[17]);
mux2 er16(i4[16],i4[0],s4,out[16]);
mux2 er17(i4[15],0,s4,out[15]);
mux2 er18(i4[14],0,s4,out[14]);
mux2 er19(i4[13],0,s4,out[13]);
mux2 er20(i4[12],0,s4,out[12]);
mux2 er21(i4[11],0,s4,out[11]);
mux2 er22(i4[10],0,s4,out[10]);
mux2 er23(i4[9],0,s4,out[9]);
mux2 er24(i4[8],0,s4,out[8]);
mux2 er25(i4[7],0,s4,out[7]);
mux2 er26(i4[6],0,s4,out[6]);
mux2 er27(i4[5],0,s4,out[5]);
mux2 er28(i4[4],0,s4,out[4]);
mux2 er29(i4[3],0,s4,out[3]);
mux2 er30(i4[2],0,s4,out[2]);
mux2 er31(i4[1],0,s4,out[1]);
mux2 er32(i4[0],0,s4,out[0]);

endmodule

module mux2(a,b,s,o);
input a,b,s;
output  o;
wire w1,w2,w3;
assign w1=~(s);
assign w2=w1&a;
assign w3=s&b;
assign o=w2|w3;
endmodule
