`include "sam.v"

module top;
reg [15:0]a,b;
reg cin,clk;
wire cout;
wire [15:0]s;

cla16 out(cout,s,a,b,cin,clk);

initial
clk=1'b0;

initial
begin


#4
a=16'b0000000000000011;
b=16'b0000000000000011;
cin=1'b1;

#4
a=16'b0000000000000011;
b=16'b0000000000000011;
cin=1'b1;


#8 $finish;
end

always
#2 clk=~clk;

initial
$monitor($time,"clock=%b,a=%b,b=%b,s=%b,cout=%b",clk,a,b,s,cout);
endmodule




