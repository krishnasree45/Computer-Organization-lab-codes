module processor(clock);


