`include "mux2.v"

module barrelshift32(a,s0,s1,s2,s3,s4,out);

input [31:0]a;
input s0,s1,s2,s3,s4;
output [31:0]out;
wire [31:0]i1,i2,i3,i4;

mux2 br1(a[31],0,s0,i1[31]);
mux2 br2(a[30],a[31],s0,i1[30]);
mux2 br3(a[29],a[30],s0,i1[29]);
mux2 br4(a[28],a[29],s0,i1[28]);
mux2 br5(a[27],a[28],s0,i1[27]);
mux2 br6(a[26],a[27],s0,i1[26]);
mux2 br7(a[25],a[26],s0,i1[25]);
mux2 br8(a[24],a[25],s0,i1[24]);
mux2 br9(a[23],a[24],s0,i1[23]);
mux2 br10(a[22],a[23],s0,i1[22]);
mux2 br11(a[21],a[22],s0,i1[21]);
mux2 br12(a[20],a[21],s0,i1[20]);
mux2 br13(a[19],a[20],s0,i1[19]);
mux2 br14(a[18],a[19],s0,i1[18]);
mux2 br15(a[17],a[18],s0,i1[17]);
mux2 br16(a[16],a[17],s0,i1[16]);
mux2 br17(a[15],a[16],s0,i1[15]);
mux2 br18(a[14],a[15],s0,i1[14]);
mux2 br19(a[13],a[14],s0,i1[13]);
mux2 br20(a[12],a[13],s0,i1[12]);
mux2 br21(a[11],a[12],s0,i1[11]);
mux2 br22(a[10],a[11],s0,i1[10]);
mux2 br23(a[9],a[10],s0,i1[9]);
mux2 br24(a[8],a[9],s0,i1[8]);
mux2 br25(a[7],a[8],s0,i1[7]);
mux2 br26(a[6],a[7],s0,i1[6]);
mux2 br27(a[5],a[6],s0,i1[5]);
mux2 br28(a[4],a[5],s0,i1[4]);
mux2 br29(a[3],a[4],s0,i1[3]);
mux2 br30(a[2],a[3],s0,i1[2]);
mux2 br31(a[1],a[2],s0,i1[1]);
mux2 br32(a[0],a[1],s0,i1[0]);


mux2 cbr1(i1[31],0,s1,i2[31]);
mux2 cbr2(i1[30],0,s1,i2[30]);
mux2 cbr3(i1[29],i1[31],s1,i2[29]);
mux2 cbr4(i1[28],i1[30],s1,i2[28]);
mux2 cbr5(i1[27],i1[29],s1,i2[27]);
mux2 cbr6(i1[26],i1[28],s1,i2[26]);
mux2 cbr7(i1[25],i1[27],s1,i2[25]);
mux2 cbr8(i1[24],i1[26],s1,i2[24]);
mux2 cbr9(i1[23],i1[25],s1,i2[23]);
mux2 cbr10(i1[22],i1[24],s1,i2[22]);
mux2 cbr11(i1[21],i1[23],s1,i2[21]);
mux2 cbr12(i1[20],i1[22],s1,i2[20]);
mux2 cbr13(i1[19],i1[21],s1,i2[19]);
mux2 cbr14(i1[18],i1[20],s1,i2[18]);
mux2 cbr15(i1[17],i1[19],s1,i2[17]);
mux2 cbr16(i1[16],i1[18],s1,i2[16]);
mux2 cbr17(i1[15],i1[17],s1,i2[15]);
mux2 cbr18(i1[14],i1[16],s1,i2[14]);
mux2 cbr19(i1[13],i1[15],s1,i2[13]);
mux2 cbr20(i1[12],i1[14],s1,i2[12]);
mux2 cbr21(i1[11],i1[13],s1,i2[11]);
mux2 cbr22(i1[10],i1[12],s1,i2[10]);
mux2 cbr23(i1[9],i1[11],s1,i2[9]);
mux2 cbr24(i1[8],i1[10],s1,i2[8]);
mux2 cbr25(i1[7],i1[9],s1,i2[7]);
mux2 cbr26(i1[6],i1[8],s1,i2[6]);
mux2 cbr27(i1[5],i1[7],s1,i2[5]);
mux2 cbr28(i1[4],i1[6],s1,i2[4]);
mux2 cbr29(i1[3],i1[5],s1,i2[3]);
mux2 cbr30(i1[2],i1[4],s1,i2[2]);
mux2 cbr31(i1[1],i1[3],s1,i2[1]);
mux2 cbr32(i1[0],i1[2],s1,i2[0]);



mux2 dbr1(i2[31],0,s2,i3[31]);
mux2 dbr2(i2[30],0,s2,i3[30]);
mux2 dbr3(i2[29],0,s2,i3[29]);
mux2 dbr4(i2[28],0,s2,i3[28]);
mux2 dbr5(i2[27],i2[31],s2,i3[27]);
mux2 dbr6(i2[26],i2[30],s2,i3[26]);
mux2 dbr7(i2[25],i2[29],s2,i3[25]);
mux2 dbr8(i2[24],i2[28],s2,i3[24]);
mux2 dbr9(i2[23],i2[27],s2,i3[23]);
mux2 dbr10(i2[22],i2[26],s2,i3[22]);
mux2 dbr11(i2[21],i2[25],s2,i3[21]);
mux2 dbr12(i2[20],i2[24],s2,i3[20]);
mux2 dbr13(i2[19],i2[23],s2,i3[19]);
mux2 dbr14(i2[18],i2[22],s2,i3[18]);
mux2 dbr15(i2[17],i2[21],s2,i3[17]);
mux2 dbr16(i2[16],i2[20],s2,i3[16]);
mux2 dbr17(i2[15],i2[19],s2,i3[15]);
mux2 dbr18(i2[14],i2[18],s2,i3[14]);
mux2 dbr19(i2[13],i2[17],s2,i3[13]);
mux2 dbr20(i2[12],i2[16],s2,i3[12]);
mux2 dbr21(i2[11],i2[15],s2,i3[11]);
mux2 dbr22(i2[10],i2[14],s2,i3[10]);
mux2 dbr23(i2[9],i2[13],s2,i3[9]);
mux2 dbr24(i2[8],i2[12],s2,i3[8]);
mux2 dbr25(i2[7],i2[11],s2,i3[7]);
mux2 dbr26(i2[6],i2[10],s2,i3[6]);
mux2 dbr27(i2[5],i2[9],s2,i3[5]);
mux2 dbr28(i2[4],i2[8],s2,i3[4]);
mux2 dbr29(i2[3],i2[7],s2,i3[3]);
mux2 dbr30(i2[2],i2[6],s2,i3[2]);
mux2 dbr31(i2[1],i2[5],s2,i3[1]);
mux2 dbr32(i2[0],i2[4],s2,i3[0]);


mux2 abr1(i3[31],0,s3,i4[31]);
mux2 abr2(i3[30],0,s3,i4[30]);
mux2 abr3(i3[29],0,s3,i4[29]);
mux2 abr4(i3[28],0,s3,i4[28]);
mux2 abr5(i3[27],0,s3,i4[27]);
mux2 abr6(i3[26],0,s3,i4[26]);
mux2 abr7(i3[25],0,s3,i4[25]);
mux2 abr8(i3[24],0,s3,i4[24]);
mux2 abr9(i3[23],i3[31],s3,i4[23]);
mux2 abr10(i3[22],i3[30],s3,i4[22]);
mux2 abr11(i3[21],i3[29],s3,i4[21]);
mux2 abr12(i3[20],i3[28],s3,i4[20]);
mux2 abr13(i3[19],i3[27],s3,i4[19]);
mux2 abr14(i3[18],i3[26],s3,i4[18]);
mux2 abr15(i3[17],i3[25],s3,i4[17]);
mux2 abr16(i3[16],i3[24],s3,i4[16]);
mux2 abr17(i3[15],i3[23],s3,i4[15]);
mux2 abr18(i3[14],i3[22],s3,i4[14]);
mux2 abr19(i3[13],i3[21],s3,i4[13]);
mux2 abr20(i3[12],i3[20],s3,i4[12]);
mux2 abr21(i3[11],i3[19],s3,i4[11]);
mux2 abr22(i3[10],i3[18],s3,i4[10]);
mux2 abr23(i3[9],i3[17],s3,i4[9]);
mux2 abr24(i3[8],i3[16],s3,i4[8]);
mux2 abr25(i3[7],i3[15],s3,i4[7]);
mux2 abr26(i3[6],i3[14],s3,i4[6]);
mux2 abr27(i3[5],i3[13],s3,i4[5]);
mux2 abr28(i3[4],i3[12],s3,i4[4]);
mux2 abr29(i3[3],i3[11],s3,i4[3]);
mux2 abr30(i3[2],i3[10],s3,i4[2]);
mux2 abr31(i3[1],i3[9],s3,i4[1]);
mux2 abr32(i3[0],i3[8],s3,i4[0]);

mux2 ebr1(i4[31],0,s4,out[31]);
mux2 ebr2(i4[30],0,s4,out[30]);
mux2 ebr3(i4[29],0,s4,out[29]);
mux2 ebr4(i4[28],0,s4,out[28]);
mux2 ebr5(i4[27],0,s4,out[27]);
mux2 ebr6(i4[26],0,s4,out[26]);
mux2 ebr7(i4[25],0,s4,out[25]);
mux2 ebr8(i4[24],0,s4,out[24]);
mux2 ebr9(i4[23],0,s4,out[23]);
mux2 ebr10(i4[22],0,s4,out[22]);
mux2 ebr11(i4[21],0,s4,out[21]);
mux2 ebr12(i4[20],0,s4,out[20]);
mux2 ebr13(i4[19],0,s4,out[19]);
mux2 ebr14(i4[18],0,s4,out[18]);
mux2 ebr15(i4[17],0,s4,out[17]);
mux2 ebr16(i4[16],0,s4,out[16]);
mux2 ebr17(i4[15],i4[31],s4,out[15]);
mux2 ebr18(i4[14],i4[30],s4,out[14]);
mux2 ebr319(i4[13],i4[29],s4,out[13]);
mux2 ebr320(i4[12],i4[28],s4,out[12]);
mux2 ebr321(i4[11],i4[27],s4,out[11]);
mux2 ebr322(i4[10],i4[26],s4,out[10]);
mux2 ebr323(i4[9],i4[25],s4,out[9]);
mux2 ebr324(i4[8],i4[24],s4,out[8]);
mux2 ebr325(i4[7],i4[23],s4,out[7]);
mux2 ebr326(i4[6],i4[22],s4,out[6]);
mux2 ebr327(i4[5],i4[21],s4,out[5]);
mux2 ebr328(i4[4],i4[20],s4,out[4]);
mux2 ebr329(i4[3],i4[19],s4,out[3]);
mux2 ebr330(i4[2],i4[18],s4,out[2]);
mux2 ebr331(i4[1],i4[17],s4,out[1]);
mux2 ebr332(i4[0],i4[16],s4,out[0]);


endmodule
