module barrellft16(a,s0,s1,s2,s3,s4,o4);
input [31:0]a;
input s0,s1,s2,s3,s4;
output [31:0]o4;
wire [31:0]o,o1,o2,o3;
wire ns0,ns1,ns2,ns3,ns4;
assign ns0=~s0;
assign ns1=~s1;
assign ns2=~s2;

assign ns3=~s3;
assign ns4=~s4;
//mux2 m33(a[31],a[32],ns0,o[32]);
mux2 m32(a[30],a[31],ns0,o[31]);
mux2 m31(a[29],a[30],ns0,o[30]);
mux2 m30(a[28],a[29],ns0,o[29]);
mux2 m29(a[27],a[28],ns0,o[28]);
mux2 m28(a[26],a[27],ns0,o[27]);
mux2 m27(a[25],a[26],ns0,o[26]);
mux2 m26(a[24],a[25],ns0,o[25]);
mux2 m25(a[23],a[24],ns0,o[24]);
mux2 m24(a[22],a[23],ns0,o[23]);
mux2 m23(a[21],a[22],ns0,o[22]);
mux2 m22(a[20],a[21],ns0,o[21]);
mux2 m21(a[19],a[20],ns0,o[20]);
mux2 m20(a[18],a[19],ns0,o[19]);
mux2 m19(a[17],a[18],ns0,o[18]);
mux2 m18(a[16],a[17],ns0,o[17]);
mux2 m17(a[15],a[16],ns0,o[16]);
mux2 m16(a[14],a[15],ns0,o[15]);
mux2 m1(a[13],a[14],ns0,o[14]);
mux2 m2(a[12],a[13],ns0,o[13]);
mux2 m3(a[11],a[12],ns0,o[12]);
mux2 m4(a[10],a[11],ns0,o[11]);
mux2 m5(a[9],a[10],ns0,o[10]);
mux2 m6(a[8],a[9],ns0,o[9]);
mux2 m7(a[7],a[8],ns0,o[8]);
mux2 m8(a[6],a[7],ns0,o[7]);
mux2 m9(a[5],a[6],ns0,o[6]);
mux2 m10(a[4],a[5],ns0,o[5]);
mux2 m11(a[3],a[4],ns0,o[4]);
mux2 m12(a[2],a[3],ns0,o[3]);
mux2 m13(a[1],a[2],ns0,o[2]);
mux2 m14(a[0],a[1],ns0,o[1]);
mux2 m15(0,a[0],ns0,o[0]);



//mux2 m33(0[30],a[32],ns0,o[32]);
mux2 M32(o[29],a[31],ns1,o1[31]);
mux2 M31(o[28],a[30],ns1,o1[30]);
mux2 M30(o[27],a[29],ns1,o1[29]);
mux2 M29(o[26],a[28],ns1,o1[28]);
mux2 M28(o[25],a[27],ns1,o1[27]);
mux2 M27(o[24],a[26],ns1,o1[26]);
mux2 M26(o[23],a[25],ns1,o1[25]);
mux2 M25(o[22],a[24],ns1,o1[24]);
mux2 M24(o[21],a[23],ns1,o1[23]);
mux2 M23(o[20],a[22],ns1,o1[22]);
mux2 M22(o[19],a[21],ns1,o1[21]);
mux2 M21(o[18],a[20],ns1,o1[20]);
mux2 M20(o[17],a[19],ns1,o1[19]);
mux2 M19(o[16],a[18],ns1,o1[18]);
mux2 M18(o[15],a[17],ns1,o1[17]);
mux2 M17(o[14],a[16],ns1,o1[16]);
mux2 M16(o[13],a[15],ns1,o1[15]);
mux2 M1(o[12],a[14],ns1,o1[14]);
mux2 M2(o[11],a[13],ns1,o1[13]);
mux2 M3(o[10],a[12],ns1,o1[12]);
mux2 M4(o[9],a[11],ns1,o1[11]);
mux2 M5(o[8],a[10],ns1,o1[10]);
mux2 M6(o[7],a[9],ns1,o1[9]);
mux2 M7(o[6],a[8],ns1,o1[8]);
mux2 M8(o[5],a[7],ns1,o1[7]);
mux2 M9(o[4],a[6],ns1,o1[6]);
mux2 M10(o[3],a[5],ns1,o1[5]);
mux2 M11(o[2],a[4],ns1,o1[4]);
mux2 M12(o[1],a[3],ns1,o1[3]);
mux2 M13(o[0],a[2],ns1,o1[2]);
mux2 M14(0,a[1],ns1,o1[1]);
mux2 M15(0,a[0],ns1,o1[0]);


mux2 R32(o1[27],o1[31],ns2,o2[31]);
mux2 R31(o1[26],o1[30],ns2,o2[30]);
mux2 R30(o1[25],o1[29],ns2,o2[29]);
mux2 R29(o1[24],o1[28],ns2,o2[28]);
mux2 R28(o1[23],o1[27],ns2,o2[27]);
mux2 R27(o1[22],o1[26],ns2,o2[26]);
mux2 R26(o1[21],o1[25],ns2,o2[25]);
mux2 R25(o1[20],o1[24],ns2,o2[24]);
mux2 R24(o1[19],o1[23],ns2,o2[23]);
mux2 R23(o1[18],o1[22],ns2,o2[22]);
mux2 R22(o1[17],o1[21],ns2,o2[21]);
mux2 R21(o1[16],o1[20],ns2,o2[20]);
mux2 R20(o1[15],o1[19],ns2,o2[19]);
mux2 R19(o1[14],o1[18],ns2,o2[18]);
mux2 R18(o1[13],o1[17],ns2,o2[17]);
mux2 R17(o1[12],o1[16],ns2,o2[16]);
mux2 R16(o1[11],o1[15],ns2,o2[15]);
mux2 R1(o1[10],o1[14],ns2,o2[14]);
mux2 R2(o1[9],o1[13],ns2,o2[13]);
mux2 R3(o1[8],o1[12],ns2,o2[12]);
mux2 R4(o1[7],o1[11],ns2,o2[11]);
mux2 R5(o1[6],o1[10],ns2,o2[10]);
mux2 R6(o1[5],o1[9],ns2,o2[9]);
mux2 R7(o1[4],o1[8],ns2,o2[8]);
mux2 R8(o1[3],o1[7],ns2,o2[7]);
mux2 R9(o1[2],o1[6],ns2,o2[6]);
mux2 R10(o1[1],o1[5],ns2,o2[5]);
mux2 R11(o1[0],o1[4],ns2,o2[4]);
mux2 R12(0,o1[3],ns2,o2[3]);
mux2 R13(0,o1[2],ns2,o2[2]);
mux2 R14(0,o1[1],ns2,o2[1]);
mux2 R15(0,o1[0],ns2,o2[0]);



mux2 S32(o2[23],o2[31],ns3,o3[31]);
mux2 S31(o2[22],o2[30],ns3,o3[30]);
mux2 S30(o2[21],o2[29],ns3,o3[29]);
mux2 S29(o2[20],o2[28],ns3,o3[28]);
mux2 S28(o2[19],o2[27],ns3,o3[27]);
mux2 S27(o2[18],o2[26],ns3,o3[26]);
mux2 S26(o2[17],o2[25],ns3,o3[25]);
mux2 S25(o2[16],o2[24],ns3,o3[24]);
mux2 S24(o2[15],o2[23],ns3,o3[23]);
mux2 S23(o2[14],o2[22],ns3,o3[22]);
mux2 S22(o2[13],o2[21],ns3,o3[21]);
mux2 S21(o2[12],o2[20],ns3,o3[20]);
mux2 S20(o2[11],o2[19],ns3,o3[19]);
mux2 S19(o2[10],o2[18],ns3,o3[18]);
mux2 S18(o2[9],o2[17],ns3,o3[17]);
mux2 S17(o2[8],o2[16],ns3,o3[16]);
mux2 S16(o2[7],o2[15],ns3,o3[15]);
mux2 S1(o2[6],o2[14],ns3,o3[14]);
mux2 S2(o2[5],o2[13],ns3,o3[13]);
mux2 S3(o2[4],o2[12],ns3,o3[12]);
mux2 S4(o2[3],o2[11],ns3,o3[11]);
mux2 S5(o2[2],o2[10],ns3,o3[10]);
mux2 S6(o2[1],o2[9],ns3,o3[9]);
mux2 S7(o2[0],o2[8],ns3,o3[8]);
mux2 S8(0,o2[7],ns3,o3[7]);
mux2 S9(0,o2[6],ns3,o3[6]);
mux2 S10(0,o2[5],ns3,o3[5]);
mux2 S11(0,o2[4],ns3,o3[4]);
mux2 S12(0,o2[3],ns3,o3[3]);
mux2 S13(0,o2[2],ns3,o3[2]);
mux2 S14(0,o2[1],ns3,o3[1]);
mux2 S15(0,o2[0],ns3,o3[0]);


mux2 L32(o3[15],o3[31],ns4,o4[31]);
mux2 L31(o3[14],o3[30],ns4,o4[30]);
mux2 L30(o3[13],o3[29],ns4,o4[29]);
mux2 L29(o3[12],o3[28],ns4,o4[28]);
mux2 L28(o3[11],o3[27],ns4,o4[27]);
mux2 L27(o3[10],o3[26],ns4,o4[26]);
mux2 L26(o3[9],o3[25],ns4,o4[25]);
mux2 L25(o3[8],o3[24],ns4,o4[24]);
mux2 L24(o3[7],o3[23],ns4,o4[23]);
mux2 L23(o3[6],o3[22],ns4,o4[22]);
mux2 L22(o3[5],o3[21],ns4,o4[21]);
mux2 L21(o3[4],o3[20],ns4,o4[20]);
mux2 L20(o3[3],o3[19],ns4,o4[19]);
mux2 L19(o3[2],o3[18],ns4,o4[18]);
mux2 L18(o3[1],o3[17],ns4,o4[17]);
mux2 L17(o3[0],o3[16],ns4,o4[16]);
mux2 L16(0,o3[15],ns4,o4[15]);
mux2 L1(0,o3[14],ns4,o4[14]);
mux2 L2(0,o3[13],ns4,o4[13]);
mux2 L3(0,o3[12],ns4,o4[12]);
mux2 L4(0,o3[11],ns4,o4[11]);
mux2 L5(0,o3[10],ns4,o4[10]);
mux2 L6(0,o3[9],ns4,o4[9]);
mux2 L7(0,o3[8],ns4,o4[8]);
mux2 L8(0,o3[7],ns4,o4[7]);
mux2 L9(0,o3[6],ns4,o4[6]);
mux2 L10(0,o3[5],ns4,o4[5]);
mux2 L11(0,o3[4],ns4,o4[4]);
mux2 L12(0,o3[3],ns4,o4[3]);
mux2 L13(0,o3[2],ns4,o4[2]);
mux2 L14(0,o3[1],ns4,o4[1]);
mux2 L15(0,o3[0],ns4,o4[0]);

endmodule

module mux2(a,b,s,o);
input a,b,s;
output  o;
wire w1,w2,w3;
assign w1=~(s);
assign w2=w1&a;
assign w3=s&b;
assign o=w2|w3;
endmodule
